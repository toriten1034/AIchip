module SystolicArray(
		input 	CLK,
		input 	RST,
		input 	WE,
		//data input
		input		[17:0]IN_0, 
		input		[17:0]IN_1, 
		input		[17:0]IN_2, 
		input		[17:0]IN_3, 
		input		[17:0]IN_4, 
		input		[17:0]IN_5, 
		input		[17:0]IN_6,
		input		[17:0]IN_7, 
		//data output 
		output	[17:0]OUT_A,
		output	[17:0]OUT_B,
		output	[17:0]OUT_C,
		output	[17:0]OUT_D,
		output	[17:0]OUT_E,
		output	[17:0]OUT_F,
		output	[17:0]OUT_G,
		output	[17:0]OUT_H

		);
	
	//row wires
	wire [17:0]A01,A12,A23,A34,A45,A56,A67;
	wire [17:0]B01,B12,B23,B34,B45,B56,B67;
	wire [17:0]C01,C12,C23,C34,C45,C56,C67;
	wire [17:0]D01,D12,D23,D34,D45,D56,D67;
	wire [17:0]E01,E12,E23,E34,E45,E56,E67;
	wire [17:0]F01,F12,F23,F34,F45,F56,F67;
	wire [17:0]G01,G12,G23,G34,G45,G56,G67;
	wire [17:0]H01,H12,H23,H34,H45,H56,H67;
	
	//col wires
	wire [17:0]AB0,AB1,AB2,AB3,AB4,AB5,AB6,AB7;
	wire [17:0]BC0,BC1,BC2,BC3,BC4,BC5,BC6,BC7;
	wire [17:0]CD0,CD1,CD2,CD3,CD4,CD5,CD6,CD7;
	wire [17:0]DE0,DE1,DE2,DE3,DE4,DE5,DE6,DE7;
	wire [17:0]EF0,EF1,EF2,EF3,EF4,EF5,EF6,EF7;
	wire [17:0]FG0,FG1,FG2,FG3,FG4,FG5,FG6,FG7;
	wire [17:0]GH0,GH1,GH2,GH3,GH4,GH5,GH6,GH7;
	
	//col 0
	PE PE_A0(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(18'b000000000_000000000),.SUMO(A01),.DIN(IN_0),.DO(AB0));
	PE PE_B0(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(18'b000000000_000000000),.SUMO(B01),.DIN(AB0), .DO(BC0));
	PE PE_C0(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(18'b000000000_000000000),.SUMO(C01),.DIN(BC0), .DO(CD0));
	PE PE_D0(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(18'b000000000_000000000),.SUMO(D01),.DIN(CD0), .DO(DE0));
	PE PE_E0(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(18'b000000000_000000000),.SUMO(E01),.DIN(DE0), .DO(EF0));
	PE PE_F0(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(18'b000000000_000000000),.SUMO(F01),.DIN(EF0), .DO(FG0));
	PE PE_G0(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(18'b000000000_000000000),.SUMO(G01),.DIN(FG0), .DO(GH0));
	PE PE_H0(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(18'b000000000_000000000),.SUMO(H01),.DIN(GH0));

	//col 1
	PE PE_A1(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(A01),.SUMO(A12),.DIN(IN_1),.DO(AB1));
	PE PE_B1(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(B01),.SUMO(B12),.DIN(AB1), .DO(BC1));
	PE PE_C1(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(C01),.SUMO(C12),.DIN(BC1), .DO(CD1));
	PE PE_D1(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(D01),.SUMO(D12),.DIN(CD1), .DO(DE1));
	PE PE_E1(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(E01),.SUMO(E12),.DIN(DE1), .DO(EF1));
	PE PE_F1(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(F01),.SUMO(F12),.DIN(EF1), .DO(FG1));
	PE PE_G1(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(G01),.SUMO(G12),.DIN(FG1), .DO(GH1));
	PE PE_H1(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(H01),.SUMO(H12),.DIN(GH1));

	//col 2
	PE PE_A2(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(A12),.SUMO(A23),.DIN(IN_2),.DO(AB2));
	PE PE_B2(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(B12),.SUMO(B23),.DIN(AB2), .DO(BC2));
	PE PE_C2(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(C12),.SUMO(C23),.DIN(BC2), .DO(CD2));
	PE PE_D2(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(D12),.SUMO(D23),.DIN(CD2), .DO(DE2));
	PE PE_E2(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(E12),.SUMO(E23),.DIN(DE2), .DO(EF2));
	PE PE_F2(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(F12),.SUMO(F23),.DIN(EF2), .DO(FG2));
	PE PE_G2(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(G12),.SUMO(G23),.DIN(FG2), .DO(GH2));
	PE PE_H2(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(H12),.SUMO(H23),.DIN(GH2));

	//col 3
	PE PE_A3(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(A23),.SUMO(A34),.DIN(IN_3),.DO(AB3));
	PE PE_B3(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(B23),.SUMO(B34),.DIN(AB3), .DO(BC3));
	PE PE_C3(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(C23),.SUMO(C34),.DIN(BC3), .DO(CD3));
	PE PE_D3(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(D23),.SUMO(D34),.DIN(CD3), .DO(DE3));
	PE PE_E3(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(E23),.SUMO(E34),.DIN(DE3), .DO(EF3));
	PE PE_F3(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(F23),.SUMO(F34),.DIN(EF3), .DO(FG3));
	PE PE_G3(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(G23),.SUMO(G34),.DIN(FG3), .DO(GH3));
	PE PE_H3(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(H23),.SUMO(H34),.DIN(GH3));

	//col 4
	PE PE_A4(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(A34),.SUMO(A45),.DIN(IN_4),.DO(AB4));
	PE PE_B4(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(B34),.SUMO(B45),.DIN(AB4), .DO(BC4));
	PE PE_C4(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(C34),.SUMO(C45),.DIN(BC4), .DO(CD4));
	PE PE_D4(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(D34),.SUMO(D45),.DIN(CD4), .DO(DE4));
	PE PE_E4(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(E34),.SUMO(E45),.DIN(DE4), .DO(EF4));
	PE PE_F4(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(F34),.SUMO(F45),.DIN(EF4), .DO(FG4));
	PE PE_G4(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(G34),.SUMO(G45),.DIN(FG4), .DO(GH4));
	PE PE_H4(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(H34),.SUMO(H45),.DIN(GH4));

	//col 5
	PE PE_A5(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(A45),.SUMO(A56),.DIN(IN_5),.DO(AB5));
	PE PE_B5(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(B45),.SUMO(B56),.DIN(AB5), .DO(BC5));
	PE PE_C5(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(C45),.SUMO(C56),.DIN(BC5), .DO(CD5));
	PE PE_D5(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(D45),.SUMO(D56),.DIN(CD5), .DO(DE5));
	PE PE_E5(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(E45),.SUMO(E56),.DIN(DE5), .DO(EF5));
	PE PE_F5(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(F45),.SUMO(F56),.DIN(EF5), .DO(FG5));
	PE PE_G5(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(G45),.SUMO(G56),.DIN(FG5), .DO(GH5));
	PE PE_H5(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(H45),.SUMO(H56),.DIN(GH5));

	//col 6
	PE PE_A6(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(A56),.SUMO(A67),.DIN(IN_6),.DO(AB6));
	PE PE_B6(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(B56),.SUMO(B67),.DIN(AB6), .DO(BC6));
	PE PE_C6(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(C56),.SUMO(C67),.DIN(BC6), .DO(CD6));
	PE PE_D6(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(D56),.SUMO(D67),.DIN(CD6), .DO(DE6));
	PE PE_E6(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(E56),.SUMO(E67),.DIN(DE6), .DO(EF6));
	PE PE_F6(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(F56),.SUMO(F67),.DIN(EF6), .DO(FG6));
	PE PE_G6(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(G56),.SUMO(G67),.DIN(FG6), .DO(GH6));
	PE PE_H6(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(H56),.SUMO(H67),.DIN(GH6));

	//col 7
	PE PE_A7(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(A67),.SUMO(OUT_A),.DIN(IN_7),.DO(AB7));
	PE PE_B7(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(B67),.SUMO(OUT_B),.DIN(AB7), .DO(BC7));
	PE PE_C7(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(C67),.SUMO(OUT_C),.DIN(BC7), .DO(CD7));
	PE PE_D7(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(D67),.SUMO(OUT_D),.DIN(CD7), .DO(DE7));
	PE PE_E7(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(E67),.SUMO(OUT_E),.DIN(DE7), .DO(EF7));
	PE PE_F7(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(F67),.SUMO(OUT_F),.DIN(EF7), .DO(FG7));
	PE PE_G7(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(G67),.SUMO(OUT_G),.DIN(FG7), .DO(GH7));
	PE PE_H7(.RST(RST),.CLK(CLK),.WE(WE),.SUMIN(H67),.SUMO(OUT_H),.DIN(GH7));

endmodule
